interface Counter_intf(input logic clk);
  logic rst;
  logic up_dn;
  logic [7:0] data_out;
  
endinterface
